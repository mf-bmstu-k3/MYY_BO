library verilog;
use verilog.vl_types.all;
entity control_unit_for_4op_BO_vlg_sample_tst is
    port(
        a               : in     vl_logic_vector(3 downto 0);
        b               : in     vl_logic_vector(3 downto 0);
        clk             : in     vl_logic;
        cop             : in     vl_logic_vector(1 downto 0);
        set             : in     vl_logic;
        sno             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end control_unit_for_4op_BO_vlg_sample_tst;
