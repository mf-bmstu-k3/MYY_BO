library verilog;
use verilog.vl_types.all;
entity alu_vhdl_vlg_vec_tst is
end alu_vhdl_vlg_vec_tst;
