library verilog;
use verilog.vl_types.all;
entity ctrl_un_BO_vlg_vec_tst is
end ctrl_un_BO_vlg_vec_tst;
