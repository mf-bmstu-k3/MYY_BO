library verilog;
use verilog.vl_types.all;
entity alu_new_vlg_vec_tst is
end alu_new_vlg_vec_tst;
