library verilog;
use verilog.vl_types.all;
entity alu_sm_vlg_vec_tst is
end alu_sm_vlg_vec_tst;
