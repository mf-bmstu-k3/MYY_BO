-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.1.0 Build 162 10/23/2013 SJ Web Edition
-- Created on Thu Nov 14 12:14:05 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SM3 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
        sno : IN STD_LOGIC := '0';
        i : IN STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
        y : OUT STD_LOGIC_VECTOR(10 DOWNTO 1);
        sko : OUT STD_LOGIC;
        incr_i : OUT STD_LOGIC
    );
END SM3;

ARCHITECTURE BEHAVIOR OF SM3 IS
    TYPE type_fstate IS (s0,s1,s2);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= s0;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,x,sno,i)
    BEGIN
        y <= "0000000000";
        sko <= '0';
        incr_i <= '0';
        CASE fstate IS
            WHEN s0 =>
                IF ((sno = '1')) THEN
                    reg_fstate <= s1;
                ELSIF (NOT((sno = '1'))) THEN
                    reg_fstate <= s0;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= s0;
                END IF;

                sko <= '0';

                IF (NOT((sno = '1'))) THEN
                    y <= "0000000000";
                ELSIF ((sno = '1')) THEN
                    y <= "0011000111";
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= "0000000000";
                END IF;
            WHEN s1 =>
                reg_fstate <= s2;

                sko <= '0';

                IF (((x(1) = '1') AND NOT((x(0) = '1')))) THEN
                    y <= "0001101000";
                ELSIF ((NOT((x(1) = '1')) AND (x(0) = '1'))) THEN
                    y <= "0001110000";
                ELSE
                    y <= "0001100000";
                END IF;
            WHEN s2 =>
                IF ((i(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= s0;
                ELSIF ((i(1 DOWNTO 0) /= "11")) THEN
                    reg_fstate <= s1;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= s2;
                END IF;

                IF ((i(1 DOWNTO 0) /= "11")) THEN
                    incr_i <= '1';
                ELSE
                    incr_i <= '0';
                END IF;

                IF ((i(1 DOWNTO 0) = "11")) THEN
                    sko <= '1';
                ELSIF ((i(1 DOWNTO 0) /= "11")) THEN
                    sko <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    sko <= '0';
                END IF;

                IF ((i(1 DOWNTO 0) /= "11")) THEN
                    y <= "0001000100";
                ELSIF ((i(1 DOWNTO 0) = "11")) THEN
                    y <= "0000000000";
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= "0000000000";
                END IF;
            WHEN OTHERS => 
                y <= "XXXXXXXXXX";
                sko <= 'X';
                incr_i <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
